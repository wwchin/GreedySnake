module red_UR_data (
	input [7:0] i_addr,
	output [23:0] head_rom_data
);
always_comb begin
		head_rom_data = {24{1'b1}};
	case(i_addr)
		0: head_rom_data = 24'h 181b1d;
		1: head_rom_data = 24'h 181b1d;
		2: head_rom_data = 24'h 181b1d;
		3: head_rom_data = 24'h cf212b;
		4: head_rom_data = 24'h f42834;
		5: head_rom_data = 24'h f42834;
		6: head_rom_data = 24'h f42834;
		7: head_rom_data = 24'h f42834;
		8: head_rom_data = 24'h f42834;
		9: head_rom_data = 24'h f42834;
		10: head_rom_data = 24'h f42834;
		11: head_rom_data = 24'h f42834;
		12: head_rom_data = 24'h cf212b;
		13: head_rom_data = 24'h 181b1d;
		14: head_rom_data = 24'h 181b1d;
		15: head_rom_data = 24'h 181b1d;
		16: head_rom_data = 24'h 181b1d;
		17: head_rom_data = 24'h 181b1d;
		18: head_rom_data = 24'h 1a1a1c;
		19: head_rom_data = 24'h cf212b;
		20: head_rom_data = 24'h f42834;
		21: head_rom_data = 24'h f42834;
		22: head_rom_data = 24'h f42834;
		23: head_rom_data = 24'h f42834;
		24: head_rom_data = 24'h f42834;
		25: head_rom_data = 24'h f42834;
		26: head_rom_data = 24'h f42834;
		27: head_rom_data = 24'h 91171f;
		28: head_rom_data = 24'h cf212b;
		29: head_rom_data = 24'h 181b1d;
		30: head_rom_data = 24'h 1a1a1c;
		31: head_rom_data = 24'h 181b1d;
		32: head_rom_data = 24'h 181b1d;
		33: head_rom_data = 24'h 181b1d;
		34: head_rom_data = 24'h 1a1a1c;
		35: head_rom_data = 24'h cf212b;
		36: head_rom_data = 24'h 91171f;
		37: head_rom_data = 24'h f42834;
		38: head_rom_data = 24'h f42834;
		39: head_rom_data = 24'h f42834;
		40: head_rom_data = 24'h f42834;
		41: head_rom_data = 24'h f42834;
		42: head_rom_data = 24'h f42834;
		43: head_rom_data = 24'h 91171f;
		44: head_rom_data = 24'h cf212b;
		45: head_rom_data = 24'h 1a1a1c;
		46: head_rom_data = 24'h 181b1d;
		47: head_rom_data = 24'h 181b1d;
		48: head_rom_data = 24'h 1a1a1c;
		49: head_rom_data = 24'h 1a1a1c;
		50: head_rom_data = 24'h 1a1a1c;
		51: head_rom_data = 24'h cf212b;
		52: head_rom_data = 24'h 91171f;
		53: head_rom_data = 24'h f42834;
		54: head_rom_data = 24'h f42834;
		55: head_rom_data = 24'h f42834;
		56: head_rom_data = 24'h f42834;
		57: head_rom_data = 24'h f42834;
		58: head_rom_data = 24'h cf212b;
		59: head_rom_data = 24'h 91171f;
		60: head_rom_data = 24'h 91171f;
		61: head_rom_data = 24'h 91171f;
		62: head_rom_data = 24'h cf212b;
		63: head_rom_data = 24'h cf212b;
		64: head_rom_data = 24'h 1a1a1c;
		65: head_rom_data = 24'h 1a1a1c;
		66: head_rom_data = 24'h 1a1a1c;
		67: head_rom_data = 24'h cf212b;
		68: head_rom_data = 24'h 91171f;
		69: head_rom_data = 24'h f42834;
		70: head_rom_data = 24'h f42834;
		71: head_rom_data = 24'h f42834;
		72: head_rom_data = 24'h f42834;
		73: head_rom_data = 24'h cf212b;
		74: head_rom_data = 24'h cf212b;
		75: head_rom_data = 24'h cf212b;
		76: head_rom_data = 24'h f42834;
		77: head_rom_data = 24'h f42834;
		78: head_rom_data = 24'h f42834;
		79: head_rom_data = 24'h f42834;
		80: head_rom_data = 24'h 1a1a1c;
		81: head_rom_data = 24'h 1a1a1c;
		82: head_rom_data = 24'h 1a1a1c;
		83: head_rom_data = 24'h cf212b;
		84: head_rom_data = 24'h 91171f;
		85: head_rom_data = 24'h f42834;
		86: head_rom_data = 24'h f42834;
		87: head_rom_data = 24'h f42834;
		88: head_rom_data = 24'h f42834;
		89: head_rom_data = 24'h cf212b;
		90: head_rom_data = 24'h cf212b;
		91: head_rom_data = 24'h f42834;
		92: head_rom_data = 24'h f42834;
		93: head_rom_data = 24'h f42834;
		94: head_rom_data = 24'h f42834;
		95: head_rom_data = 24'h f42834;
		96: head_rom_data = 24'h 1a1a1c;
		97: head_rom_data = 24'h 1a1a1c;
		98: head_rom_data = 24'h 1a1a1c;
		99: head_rom_data = 24'h cf212b;
		100: head_rom_data = 24'h f42834;
		101: head_rom_data = 24'h f42834;
		102: head_rom_data = 24'h f42834;
		103: head_rom_data = 24'h f42834;
		104: head_rom_data = 24'h f42834;
		105: head_rom_data = 24'h f42834;
		106: head_rom_data = 24'h f42834;
		107: head_rom_data = 24'h f42834;
		108: head_rom_data = 24'h f42834;
		109: head_rom_data = 24'h f42834;
		110: head_rom_data = 24'h f42834;
		111: head_rom_data = 24'h f42834;
		112: head_rom_data = 24'h 1a1a1c;
		113: head_rom_data = 24'h 1a1a1c;
		114: head_rom_data = 24'h 1a1a1c;
		115: head_rom_data = 24'h cf212b;
		116: head_rom_data = 24'h f42834;
		117: head_rom_data = 24'h f42834;
		118: head_rom_data = 24'h f42834;
		119: head_rom_data = 24'h cf212b;
		120: head_rom_data = 24'h cf212b;
		121: head_rom_data = 24'h f42834;
		122: head_rom_data = 24'h f42834;
		123: head_rom_data = 24'h f42834;
		124: head_rom_data = 24'h f42834;
		125: head_rom_data = 24'h f42834;
		126: head_rom_data = 24'h f42834;
		127: head_rom_data = 24'h f42834;
		128: head_rom_data = 24'h 1a1a1c;
		129: head_rom_data = 24'h 1a1a1c;
		130: head_rom_data = 24'h 1a1a1c;
		131: head_rom_data = 24'h cf212b;
		132: head_rom_data = 24'h cf212b;
		133: head_rom_data = 24'h 91171f;
		134: head_rom_data = 24'h cf212b;
		135: head_rom_data = 24'h cf212b;
		136: head_rom_data = 24'h cf212b;
		137: head_rom_data = 24'h f42834;
		138: head_rom_data = 24'h f42834;
		139: head_rom_data = 24'h f42834;
		140: head_rom_data = 24'h f42834;
		141: head_rom_data = 24'h f42834;
		142: head_rom_data = 24'h f42834;
		143: head_rom_data = 24'h f42834;
		144: head_rom_data = 24'h 1a1a1c;
		145: head_rom_data = 24'h 1a1a1c;
		146: head_rom_data = 24'h 1a1a1c;
		147: head_rom_data = 24'h 1a1a1c;
		148: head_rom_data = 24'h cf212b;
		149: head_rom_data = 24'h 91171f;
		150: head_rom_data = 24'h 91171f;
		151: head_rom_data = 24'h cf212b;
		152: head_rom_data = 24'h f42834;
		153: head_rom_data = 24'h f42834;
		154: head_rom_data = 24'h f42834;
		155: head_rom_data = 24'h f42834;
		156: head_rom_data = 24'h f42834;
		157: head_rom_data = 24'h f42834;
		158: head_rom_data = 24'h f42834;
		159: head_rom_data = 24'h f42834;
		160: head_rom_data = 24'h 1a1a1c;
		161: head_rom_data = 24'h 1a1a1c;
		162: head_rom_data = 24'h 1a1a1c;
		163: head_rom_data = 24'h 1a1a1c;
		164: head_rom_data = 24'h 1a1a1c;
		165: head_rom_data = 24'h cf212b;
		166: head_rom_data = 24'h 91171f;
		167: head_rom_data = 24'h 91171f;
		168: head_rom_data = 24'h f42834;
		169: head_rom_data = 24'h f42834;
		170: head_rom_data = 24'h f42834;
		171: head_rom_data = 24'h f42834;
		172: head_rom_data = 24'h f42834;
		173: head_rom_data = 24'h f42834;
		174: head_rom_data = 24'h f42834;
		175: head_rom_data = 24'h f42834;
		176: head_rom_data = 24'h 1a1a1c;
		177: head_rom_data = 24'h 1a1a1c;
		178: head_rom_data = 24'h 1a1a1c;
		179: head_rom_data = 24'h 1a1a1c;
		180: head_rom_data = 24'h 1a1a1c;
		181: head_rom_data = 24'h 1a1a1c;
		182: head_rom_data = 24'h cf212b;
		183: head_rom_data = 24'h 91171f;
		184: head_rom_data = 24'h f42834;
		185: head_rom_data = 24'h f42834;
		186: head_rom_data = 24'h f42834;
		187: head_rom_data = 24'h f42834;
		188: head_rom_data = 24'h f42834;
		189: head_rom_data = 24'h f42834;
		190: head_rom_data = 24'h f42834;
		191: head_rom_data = 24'h f42834;
		192: head_rom_data = 24'h 1a1a1c;
		193: head_rom_data = 24'h 1a1a1c;
		194: head_rom_data = 24'h 1a1a1c;
		195: head_rom_data = 24'h 1a1a1c;
		196: head_rom_data = 24'h 1a1a1c;
		197: head_rom_data = 24'h 1a1a1c;
		198: head_rom_data = 24'h cf212b;
		199: head_rom_data = 24'h cf212b;
		200: head_rom_data = 24'h cf212b;
		201: head_rom_data = 24'h cf212b;
		202: head_rom_data = 24'h 91171f;
		203: head_rom_data = 24'h 91171f;
		204: head_rom_data = 24'h 91171f;
		205: head_rom_data = 24'h 91171f;
		206: head_rom_data = 24'h cf212b;
		207: head_rom_data = 24'h cf212b;
		208: head_rom_data = 24'h 1a1a1c;
		209: head_rom_data = 24'h 1a1a1c;
		210: head_rom_data = 24'h 1a1a1c;
		211: head_rom_data = 24'h 1a1a1c;
		212: head_rom_data = 24'h 1a1a1c;
		213: head_rom_data = 24'h 1a1a1c;
		214: head_rom_data = 24'h 1a1a1c;
		215: head_rom_data = 24'h 1a1a1c;
		216: head_rom_data = 24'h 1a1a1c;
		217: head_rom_data = 24'h 1a1a1c;
		218: head_rom_data = 24'h 1a1a1c;
		219: head_rom_data = 24'h 1a1a1c;
		220: head_rom_data = 24'h 1a1a1c;
		221: head_rom_data = 24'h 1a1a1c;
		222: head_rom_data = 24'h 1a1a1c;
		223: head_rom_data = 24'h 181b1d;
		224: head_rom_data = 24'h 1a1a1c;
		225: head_rom_data = 24'h 1a1a1c;
		226: head_rom_data = 24'h 1a1a1c;
		227: head_rom_data = 24'h 1a1a1c;
		228: head_rom_data = 24'h 181b1d;
		229: head_rom_data = 24'h 181b1d;
		230: head_rom_data = 24'h 181b1d;
		231: head_rom_data = 24'h 181b1d;
		232: head_rom_data = 24'h 181b1d;
		233: head_rom_data = 24'h 181b1d;
		234: head_rom_data = 24'h 181b1d;
		235: head_rom_data = 24'h 181b1d;
		236: head_rom_data = 24'h 181b1d;
		237: head_rom_data = 24'h 181b1d;
		238: head_rom_data = 24'h 181b1d;
		239: head_rom_data = 24'h 181b1d;
		240: head_rom_data = 24'h 1a1a1c;
		241: head_rom_data = 24'h 1a1a1c;
		242: head_rom_data = 24'h 1a1a1c;
		243: head_rom_data = 24'h 1a1a1c;
		244: head_rom_data = 24'h 181b1d;
		245: head_rom_data = 24'h 181b1d;
		246: head_rom_data = 24'h 181b1d;
		247: head_rom_data = 24'h 181b1d;
		248: head_rom_data = 24'h 181b1d;
		249: head_rom_data = 24'h 181b1d;
		250: head_rom_data = 24'h 181b1d;
		251: head_rom_data = 24'h 181b1d;
		252: head_rom_data = 24'h 181b1d;
		253: head_rom_data = 24'h 181b1d;
		254: head_rom_data = 24'h 181b1d;
		255: head_rom_data = 24'h 181b1d;
		default: ;
	endcase
end

endmodule