module green_tail_data (
	input [7:0] i_addr,
	output [23:0] head_rom_data
);
always_comb begin
	case(i_addr)
		0: head_rom_data = 24'h 181b1d;
		1: head_rom_data = 24'h 181b1d;
		2: head_rom_data = 24'h 181b1d;
		3: head_rom_data = 24'h 074b2b;
		4: head_rom_data = 24'h c3ed80;
		5: head_rom_data = 24'h c3ed80;
		6: head_rom_data = 24'h c3ed80;
		7: head_rom_data = 24'h c3ed80;
		8: head_rom_data = 24'h c3ed80;
		9: head_rom_data = 24'h c3ed80;
		10: head_rom_data = 24'h c3ed80;
		11: head_rom_data = 24'h c3ed80;
		12: head_rom_data = 24'h 074b2b;
		13: head_rom_data = 24'h 181b1d;
		14: head_rom_data = 24'h 181b1d;
		15: head_rom_data = 24'h 181b1d;
		16: head_rom_data = 24'h 181b1d;
		17: head_rom_data = 24'h 181b1d;
		18: head_rom_data = 24'h 181b1d;
		19: head_rom_data = 24'h 074b2b;
		20: head_rom_data = 24'h c3ed80;
		21: head_rom_data = 24'h c3ed80;
		22: head_rom_data = 24'h c3ed80;
		23: head_rom_data = 24'h c3ed80;
		24: head_rom_data = 24'h c3ed80;
		25: head_rom_data = 24'h c3ed80;
		26: head_rom_data = 24'h c3ed80;
		27: head_rom_data = 24'h c3ed80;
		28: head_rom_data = 24'h 074b2b;
		29: head_rom_data = 24'h 181b1d;
		30: head_rom_data = 24'h 181b1d;
		31: head_rom_data = 24'h 181b1d;
		32: head_rom_data = 24'h 181b1d;
		33: head_rom_data = 24'h 181b1d;
		34: head_rom_data = 24'h 181b1d;
		35: head_rom_data = 24'h 074b2b;
		36: head_rom_data = 24'h c3ed80;
		37: head_rom_data = 24'h c3ed80;
		38: head_rom_data = 24'h c3ed80;
		39: head_rom_data = 24'h c3ed80;
		40: head_rom_data = 24'h c3ed80;
		41: head_rom_data = 24'h c3ed80;
		42: head_rom_data = 24'h c3ed80;
		43: head_rom_data = 24'h c3ed80;
		44: head_rom_data = 24'h 074b2b;
		45: head_rom_data = 24'h 181b1d;
		46: head_rom_data = 24'h 181b1d;
		47: head_rom_data = 24'h 181b1d;
		48: head_rom_data = 24'h 181b1d;
		49: head_rom_data = 24'h 181b1d;
		50: head_rom_data = 24'h 181b1d;
		51: head_rom_data = 24'h 074b2b;
		52: head_rom_data = 24'h 85bf2f;
		53: head_rom_data = 24'h 85bf2f;
		54: head_rom_data = 24'h 85bf2f;
		55: head_rom_data = 24'h c3ed80;
		56: head_rom_data = 24'h c3ed80;
		57: head_rom_data = 24'h 85bf2f;
		58: head_rom_data = 24'h 85bf2f;
		59: head_rom_data = 24'h 85bf2f;
		60: head_rom_data = 24'h 074b2b;
		61: head_rom_data = 24'h 181b1d;
		62: head_rom_data = 24'h 181b1d;
		63: head_rom_data = 24'h 181b1d;
		64: head_rom_data = 24'h 181b1d;
		65: head_rom_data = 24'h 181b1d;
		66: head_rom_data = 24'h 181b1d;
		67: head_rom_data = 24'h 074b2b;
		68: head_rom_data = 24'h 85bf2f;
		69: head_rom_data = 24'h 85bf2f;
		70: head_rom_data = 24'h 85bf2f;
		71: head_rom_data = 24'h c3ed80;
		72: head_rom_data = 24'h c3ed80;
		73: head_rom_data = 24'h 85bf2f;
		74: head_rom_data = 24'h 85bf2f;
		75: head_rom_data = 24'h 85bf2f;
		76: head_rom_data = 24'h 074b2b;
		77: head_rom_data = 24'h 181b1d;
		78: head_rom_data = 24'h 181b1d;
		79: head_rom_data = 24'h 181b1d;
		80: head_rom_data = 24'h 181b1d;
		81: head_rom_data = 24'h 181b1d;
		82: head_rom_data = 24'h 181b1d;
		83: head_rom_data = 24'h 074b2b;
		84: head_rom_data = 24'h c3ed80;
		85: head_rom_data = 24'h c3ed80;
		86: head_rom_data = 24'h c3ed80;
		87: head_rom_data = 24'h c3ed80;
		88: head_rom_data = 24'h c3ed80;
		89: head_rom_data = 24'h c3ed80;
		90: head_rom_data = 24'h c3ed80;
		91: head_rom_data = 24'h c3ed80;
		92: head_rom_data = 24'h 074b2b;
		93: head_rom_data = 24'h 181b1d;
		94: head_rom_data = 24'h 181b1d;
		95: head_rom_data = 24'h 181b1d;
		96: head_rom_data = 24'h 181b1d;
		97: head_rom_data = 24'h 181b1d;
		98: head_rom_data = 24'h 181b1d;
		99: head_rom_data = 24'h 074b2b;
		100: head_rom_data = 24'h c3ed80;
		101: head_rom_data = 24'h c3ed80;
		102: head_rom_data = 24'h c3ed80;
		103: head_rom_data = 24'h c3ed80;
		104: head_rom_data = 24'h c3ed80;
		105: head_rom_data = 24'h c3ed80;
		106: head_rom_data = 24'h c3ed80;
		107: head_rom_data = 24'h c3ed80;
		108: head_rom_data = 24'h 074b2b;
		109: head_rom_data = 24'h 181b1d;
		110: head_rom_data = 24'h 181b1d;
		111: head_rom_data = 24'h 181b1d;
		112: head_rom_data = 24'h 181b1d;
		113: head_rom_data = 24'h 181b1d;
		114: head_rom_data = 24'h 181b1d;
		115: head_rom_data = 24'h 074b2b;
		116: head_rom_data = 24'h c3ed80;
		117: head_rom_data = 24'h c3ed80;
		118: head_rom_data = 24'h c3ed80;
		119: head_rom_data = 24'h 9ce238;
		120: head_rom_data = 24'h 9ce238;
		121: head_rom_data = 24'h c3ed80;
		122: head_rom_data = 24'h c3ed80;
		123: head_rom_data = 24'h c3ed80;
		124: head_rom_data = 24'h 074b2b;
		125: head_rom_data = 24'h 181b1d;
		126: head_rom_data = 24'h 181b1d;
		127: head_rom_data = 24'h 181b1d;
		128: head_rom_data = 24'h 181b1d;
		129: head_rom_data = 24'h 181b1d;
		130: head_rom_data = 24'h 181b1d;
		131: head_rom_data = 24'h 074b2b;
		132: head_rom_data = 24'h 5d8721;
		133: head_rom_data = 24'h c3ed80;
		134: head_rom_data = 24'h c3ed80;
		135: head_rom_data = 24'h 9ce238;
		136: head_rom_data = 24'h 9ce238;
		137: head_rom_data = 24'h c3ed80;
		138: head_rom_data = 24'h c3ed80;
		139: head_rom_data = 24'h 5d8721;
		140: head_rom_data = 24'h 074b2b;
		141: head_rom_data = 24'h 181b1d;
		142: head_rom_data = 24'h 181b1d;
		143: head_rom_data = 24'h 181b1d;
		144: head_rom_data = 24'h 181b1d;
		145: head_rom_data = 24'h 181b1d;
		146: head_rom_data = 24'h 181b1d;
		147: head_rom_data = 24'h 074b2b;
		148: head_rom_data = 24'h 5d8721;
		149: head_rom_data = 24'h c3ed80;
		150: head_rom_data = 24'h c3ed80;
		151: head_rom_data = 24'h c3ed80;
		152: head_rom_data = 24'h c3ed80;
		153: head_rom_data = 24'h c3ed80;
		154: head_rom_data = 24'h c3ed80;
		155: head_rom_data = 24'h 5d8721;
		156: head_rom_data = 24'h 074b2b;
		157: head_rom_data = 24'h 181b1d;
		158: head_rom_data = 24'h 181b1d;
		159: head_rom_data = 24'h 181b1d;
		160: head_rom_data = 24'h 181b1d;
		161: head_rom_data = 24'h 181b1d;
		162: head_rom_data = 24'h 181b1d;
		163: head_rom_data = 24'h 181b1d;
		164: head_rom_data = 24'h 074b2b;
		165: head_rom_data = 24'h c3ed80;
		166: head_rom_data = 24'h c3ed80;
		167: head_rom_data = 24'h c3ed80;
		168: head_rom_data = 24'h c3ed80;
		169: head_rom_data = 24'h c3ed80;
		170: head_rom_data = 24'h c3ed80;
		171: head_rom_data = 24'h 074b2b;
		172: head_rom_data = 24'h 181b1d;
		173: head_rom_data = 24'h 181b1d;
		174: head_rom_data = 24'h 181b1d;
		175: head_rom_data = 24'h 181b1d;
		176: head_rom_data = 24'h 181b1d;
		177: head_rom_data = 24'h 181b1d;
		178: head_rom_data = 24'h 181b1d;
		179: head_rom_data = 24'h 181b1d;
		180: head_rom_data = 24'h 074b2b;
		181: head_rom_data = 24'h 5d8721;
		182: head_rom_data = 24'h 5d8721;
		183: head_rom_data = 24'h c3ed80;
		184: head_rom_data = 24'h c3ed80;
		185: head_rom_data = 24'h 5d8721;
		186: head_rom_data = 24'h 5d8721;
		187: head_rom_data = 24'h 074b2b;
		188: head_rom_data = 24'h 181b1d;
		189: head_rom_data = 24'h 181b1d;
		190: head_rom_data = 24'h 181b1d;
		191: head_rom_data = 24'h 181b1d;
		192: head_rom_data = 24'h 181b1d;
		193: head_rom_data = 24'h 181b1d;
		194: head_rom_data = 24'h 181b1d;
		195: head_rom_data = 24'h 181b1d;
		196: head_rom_data = 24'h 074b2b;
		197: head_rom_data = 24'h 074b2b;
		198: head_rom_data = 24'h 5d8721;
		199: head_rom_data = 24'h c3ed80;
		200: head_rom_data = 24'h c3ed80;
		201: head_rom_data = 24'h 5d8721;
		202: head_rom_data = 24'h 074b2b;
		203: head_rom_data = 24'h 074b2b;
		204: head_rom_data = 24'h 181b1d;
		205: head_rom_data = 24'h 181b1d;
		206: head_rom_data = 24'h 181b1d;
		207: head_rom_data = 24'h 181b1d;
		208: head_rom_data = 24'h 181b1d;
		209: head_rom_data = 24'h 181b1d;
		210: head_rom_data = 24'h 181b1d;
		211: head_rom_data = 24'h 181b1d;
		212: head_rom_data = 24'h 181b1d;
		213: head_rom_data = 24'h 181b1d;
		214: head_rom_data = 24'h 074b2b;
		215: head_rom_data = 24'h c3ed80;
		216: head_rom_data = 24'h c3ed80;
		217: head_rom_data = 24'h 074b2b;
		218: head_rom_data = 24'h 181b1d;
		219: head_rom_data = 24'h 181b1d;
		220: head_rom_data = 24'h 181b1d;
		221: head_rom_data = 24'h 181b1d;
		222: head_rom_data = 24'h 181b1d;
		223: head_rom_data = 24'h 181b1d;
		224: head_rom_data = 24'h 181b1d;
		225: head_rom_data = 24'h 181b1d;
		226: head_rom_data = 24'h 181b1d;
		227: head_rom_data = 24'h 181b1d;
		228: head_rom_data = 24'h 181b1d;
		229: head_rom_data = 24'h 181b1d;
		230: head_rom_data = 24'h 074b2b;
		231: head_rom_data = 24'h 5d8721;
		232: head_rom_data = 24'h 5d8721;
		233: head_rom_data = 24'h 074b2b;
		234: head_rom_data = 24'h 181b1d;
		235: head_rom_data = 24'h 181b1d;
		236: head_rom_data = 24'h 181b1d;
		237: head_rom_data = 24'h 181b1d;
		238: head_rom_data = 24'h 181b1d;
		239: head_rom_data = 24'h 181b1d;
		240: head_rom_data = 24'h 181b1d;
		241: head_rom_data = 24'h 181b1d;
		242: head_rom_data = 24'h 181b1d;
		243: head_rom_data = 24'h 181b1d;
		244: head_rom_data = 24'h 181b1d;
		245: head_rom_data = 24'h 181b1d;
		246: head_rom_data = 24'h 181b1d;
		247: head_rom_data = 24'h 07443a;
		248: head_rom_data = 24'h 07443a;
		249: head_rom_data = 24'h 181b1d;
		250: head_rom_data = 24'h 181b1d;
		251: head_rom_data = 24'h 181b1d;
		252: head_rom_data = 24'h 181b1d;
		253: head_rom_data = 24'h 181b1d;
		254: head_rom_data = 24'h 181b1d;
		255: head_rom_data = 24'h 181b1d;
		default: ;
	endcase
end

endmodule