module green_head_data (
	input [7:0] i_addr,
	output [23:0] head_rom_data
);
always_comb begin
	case(i_addr)
		0: head_rom_data = 24'h 1a1a1c;
		1: head_rom_data = 24'h 1a1a1c;
		2: head_rom_data = 24'h 1a1a1c;
		3: head_rom_data = 24'h 1a1a1c;
		4: head_rom_data = 24'h 1a1a1c;
		5: head_rom_data = 24'h cf212b;
		6: head_rom_data = 24'h 1a1a1c;
		7: head_rom_data = 24'h 1a1a1c;
		8: head_rom_data = 24'h 1a1a1c;
		9: head_rom_data = 24'h 1a1a1c;
		10: head_rom_data = 24'h cf212b;
		11: head_rom_data = 24'h 1a1a1c;
		12: head_rom_data = 24'h 1a1a1c;
		13: head_rom_data = 24'h 1a1a1c;
		14: head_rom_data = 24'h 1a1a1c;
		15: head_rom_data = 24'h 1a1a1c;
		16: head_rom_data = 24'h 1a1a1c;
		17: head_rom_data = 24'h 1a1a1c;
		18: head_rom_data = 24'h 1a1a1c;
		19: head_rom_data = 24'h 1a1a1c;
		20: head_rom_data = 24'h 1a1a1c;
		21: head_rom_data = 24'h 1a1a1c;
		22: head_rom_data = 24'h cf212b;
		23: head_rom_data = 24'h 1a1a1c;
		24: head_rom_data = 24'h 1a1a1c;
		25: head_rom_data = 24'h cf212b;
		26: head_rom_data = 24'h 1a1a1c;
		27: head_rom_data = 24'h 1a1a1c;
		28: head_rom_data = 24'h 1a1a1c;
		29: head_rom_data = 24'h 1a1a1c;
		30: head_rom_data = 24'h 1a1a1c;
		31: head_rom_data = 24'h 1a1a1c;
		32: head_rom_data = 24'h 1a1a1c;
		33: head_rom_data = 24'h 1a1a1c;
		34: head_rom_data = 24'h 1a1a1c;
		35: head_rom_data = 24'h 1a1a1c;
		36: head_rom_data = 24'h 1a1a1c;
		37: head_rom_data = 24'h 1a1a1c;
		38: head_rom_data = 24'h 181b1d;
		39: head_rom_data = 24'h cf212b;
		40: head_rom_data = 24'h cf212b;
		41: head_rom_data = 24'h 181b1d;
		42: head_rom_data = 24'h 1a1a1c;
		43: head_rom_data = 24'h 1a1a1c;
		44: head_rom_data = 24'h 1a1a1c;
		45: head_rom_data = 24'h 1a1a1c;
		46: head_rom_data = 24'h 1a1a1c;
		47: head_rom_data = 24'h 1a1a1c;
		48: head_rom_data = 24'h 1a1a1c;
		49: head_rom_data = 24'h 1a1a1c;
		50: head_rom_data = 24'h 1a1a1c;
		51: head_rom_data = 24'h 1a1a1c;
		52: head_rom_data = 24'h 074b2b;
		53: head_rom_data = 24'h 074b2b;
		54: head_rom_data = 24'h 074b2b;
		55: head_rom_data = 24'h cf212b;
		56: head_rom_data = 24'h cf212b;
		57: head_rom_data = 24'h 074b2b;
		58: head_rom_data = 24'h 074b2b;
		59: head_rom_data = 24'h 074b2b;
		60: head_rom_data = 24'h 1a1a1c;
		61: head_rom_data = 24'h 1a1a1c;
		62: head_rom_data = 24'h 1a1a1c;
		63: head_rom_data = 24'h 1a1a1c;
		64: head_rom_data = 24'h 1a1a1c;
		65: head_rom_data = 24'h 1a1a1c;
		66: head_rom_data = 24'h 1a1a1c;
		67: head_rom_data = 24'h 1a1a1c;
		68: head_rom_data = 24'h 074b2b;
		69: head_rom_data = 24'h c3ed80;
		70: head_rom_data = 24'h c3ed80;
		71: head_rom_data = 24'h cf212b;
		72: head_rom_data = 24'h cf212b;
		73: head_rom_data = 24'h c3ed80;
		74: head_rom_data = 24'h c3ed80;
		75: head_rom_data = 24'h 074b2b;
		76: head_rom_data = 24'h 1a1a1c;
		77: head_rom_data = 24'h 1a1a1c;
		78: head_rom_data = 24'h 1a1a1c;
		79: head_rom_data = 24'h 1a1a1c;
		80: head_rom_data = 24'h 1a1a1c;
		81: head_rom_data = 24'h 1a1a1c;
		82: head_rom_data = 24'h 1a1a1c;
		83: head_rom_data = 24'h 074b2b;
		84: head_rom_data = 24'h 074b2b;
		85: head_rom_data = 24'h c3ed80;
		86: head_rom_data = 24'h c3ed80;
		87: head_rom_data = 24'h c3ed80;
		88: head_rom_data = 24'h c3ed80;
		89: head_rom_data = 24'h c3ed80;
		90: head_rom_data = 24'h c3ed80;
		91: head_rom_data = 24'h 074b2b;
		92: head_rom_data = 24'h 074b2b;
		93: head_rom_data = 24'h 1a1a1c;
		94: head_rom_data = 24'h 1a1a1c;
		95: head_rom_data = 24'h 1a1a1c;
		96: head_rom_data = 24'h 1a1a1c;
		97: head_rom_data = 24'h 1a1a1c;
		98: head_rom_data = 24'h 1a1a1c;
		99: head_rom_data = 24'h 074b2b;
		100: head_rom_data = 24'h c3ed80;
		101: head_rom_data = 24'h c3ed80;
		102: head_rom_data = 24'h c3ed80;
		103: head_rom_data = 24'h c3ed80;
		104: head_rom_data = 24'h c3ed80;
		105: head_rom_data = 24'h c3ed80;
		106: head_rom_data = 24'h c3ed80;
		107: head_rom_data = 24'h c3ed80;
		108: head_rom_data = 24'h 074b2b;
		109: head_rom_data = 24'h 1a1a1c;
		110: head_rom_data = 24'h 1a1a1c;
		111: head_rom_data = 24'h 1a1a1c;
		112: head_rom_data = 24'h 1a1a1c;
		113: head_rom_data = 24'h 1a1a1c;
		114: head_rom_data = 24'h 1a1a1c;
		115: head_rom_data = 24'h 074b2b;
		116: head_rom_data = 24'h c3ed80;
		117: head_rom_data = 24'h 1a1a1c;
		118: head_rom_data = 24'h ffffff;
		119: head_rom_data = 24'h c3ed80;
		120: head_rom_data = 24'h c3ed80;
		121: head_rom_data = 24'h ffffff;
		122: head_rom_data = 24'h 1a1a1c;
		123: head_rom_data = 24'h c3ed80;
		124: head_rom_data = 24'h 074b2b;
		125: head_rom_data = 24'h 1a1a1c;
		126: head_rom_data = 24'h 1a1a1c;
		127: head_rom_data = 24'h 1a1a1c;
		128: head_rom_data = 24'h 1a1a1c;
		129: head_rom_data = 24'h 1a1a1c;
		130: head_rom_data = 24'h 1a1a1c;
		131: head_rom_data = 24'h 074b2b;
		132: head_rom_data = 24'h c3ed80;
		133: head_rom_data = 24'h 1a1a1c;
		134: head_rom_data = 24'h 1a1a1c;
		135: head_rom_data = 24'h c3ed80;
		136: head_rom_data = 24'h c3ed80;
		137: head_rom_data = 24'h 1a1a1c;
		138: head_rom_data = 24'h 1a1a1c;
		139: head_rom_data = 24'h c3ed80;
		140: head_rom_data = 24'h 074b2b;
		141: head_rom_data = 24'h 1a1a1c;
		142: head_rom_data = 24'h 1a1a1c;
		143: head_rom_data = 24'h 1a1a1c;
		144: head_rom_data = 24'h 1a1a1c;
		145: head_rom_data = 24'h 1a1a1c;
		146: head_rom_data = 24'h 1a1a1c;
		147: head_rom_data = 24'h 074b2b;
		148: head_rom_data = 24'h c3ed80;
		149: head_rom_data = 24'h c3ed80;
		150: head_rom_data = 24'h c3ed80;
		151: head_rom_data = 24'h c3ed80;
		152: head_rom_data = 24'h c3ed80;
		153: head_rom_data = 24'h c3ed80;
		154: head_rom_data = 24'h c3ed80;
		155: head_rom_data = 24'h c3ed80;
		156: head_rom_data = 24'h 074b2b;
		157: head_rom_data = 24'h 1a1a1c;
		158: head_rom_data = 24'h 1a1a1c;
		159: head_rom_data = 24'h 1a1a1c;
		160: head_rom_data = 24'h 1a1a1c;
		161: head_rom_data = 24'h 1a1a1c;
		162: head_rom_data = 24'h 1a1a1c;
		163: head_rom_data = 24'h 074b2b;
		164: head_rom_data = 24'h c3ed80;
		165: head_rom_data = 24'h c3ed80;
		166: head_rom_data = 24'h c3ed80;
		167: head_rom_data = 24'h 85bf2f;
		168: head_rom_data = 24'h 85bf2f;
		169: head_rom_data = 24'h c3ed80;
		170: head_rom_data = 24'h c3ed80;
		171: head_rom_data = 24'h c3ed80;
		172: head_rom_data = 24'h 074b2b;
		173: head_rom_data = 24'h 1a1a1c;
		174: head_rom_data = 24'h 1a1a1c;
		175: head_rom_data = 24'h 1a1a1c;
		176: head_rom_data = 24'h 1a1a1c;
		177: head_rom_data = 24'h 1a1a1c;
		178: head_rom_data = 24'h 1a1a1c;
		179: head_rom_data = 24'h 074b2b;
		180: head_rom_data = 24'h 5d8721;
		181: head_rom_data = 24'h c3ed80;
		182: head_rom_data = 24'h c3ed80;
		183: head_rom_data = 24'h c3ed80;
		184: head_rom_data = 24'h c3ed80;
		185: head_rom_data = 24'h c3ed80;
		186: head_rom_data = 24'h c3ed80;
		187: head_rom_data = 24'h 5d8721;
		188: head_rom_data = 24'h 074b2b;
		189: head_rom_data = 24'h 1a1a1c;
		190: head_rom_data = 24'h 1a1a1c;
		191: head_rom_data = 24'h 1a1a1c;
		192: head_rom_data = 24'h 1a1a1c;
		193: head_rom_data = 24'h 1a1a1c;
		194: head_rom_data = 24'h 1a1a1c;
		195: head_rom_data = 24'h 074b2b;
		196: head_rom_data = 24'h 5d8721;
		197: head_rom_data = 24'h c3ed80;
		198: head_rom_data = 24'h c3ed80;
		199: head_rom_data = 24'h c3ed80;
		200: head_rom_data = 24'h c3ed80;
		201: head_rom_data = 24'h c3ed80;
		202: head_rom_data = 24'h c3ed80;
		203: head_rom_data = 24'h 5d8721;
		204: head_rom_data = 24'h 074b2b;
		205: head_rom_data = 24'h 1a1a1c;
		206: head_rom_data = 24'h 1a1a1c;
		207: head_rom_data = 24'h 1a1a1c;
		208: head_rom_data = 24'h 1a1a1c;
		209: head_rom_data = 24'h 1a1a1c;
		210: head_rom_data = 24'h 1a1a1c;
		211: head_rom_data = 24'h 074b2b;
		212: head_rom_data = 24'h c3ed80;
		213: head_rom_data = 24'h c3ed80;
		214: head_rom_data = 24'h 85bf2f;
		215: head_rom_data = 24'h 85bf2f;
		216: head_rom_data = 24'h 85bf2f;
		217: head_rom_data = 24'h 85bf2f;
		218: head_rom_data = 24'h c3ed80;
		219: head_rom_data = 24'h c3ed80;
		220: head_rom_data = 24'h 074b2b;
		221: head_rom_data = 24'h 1a1a1c;
		222: head_rom_data = 24'h 1a1a1c;
		223: head_rom_data = 24'h 1a1a1c;
		224: head_rom_data = 24'h 1a1a1c;
		225: head_rom_data = 24'h 1a1a1c;
		226: head_rom_data = 24'h 1a1a1c;
		227: head_rom_data = 24'h 074b2b;
		228: head_rom_data = 24'h c3ed80;
		229: head_rom_data = 24'h c3ed80;
		230: head_rom_data = 24'h 85bf2f;
		231: head_rom_data = 24'h 85bf2f;
		232: head_rom_data = 24'h 85bf2f;
		233: head_rom_data = 24'h 85bf2f;
		234: head_rom_data = 24'h c3ed80;
		235: head_rom_data = 24'h c3ed80;
		236: head_rom_data = 24'h 074b2b;
		237: head_rom_data = 24'h 1a1a1c;
		238: head_rom_data = 24'h 1a1a1c;
		239: head_rom_data = 24'h 1a1a1c;
		240: head_rom_data = 24'h 1a1a1c;
		241: head_rom_data = 24'h 1a1a1c;
		242: head_rom_data = 24'h 1a1a1c;
		243: head_rom_data = 24'h 074b2b;
		244: head_rom_data = 24'h c3ed80;
		245: head_rom_data = 24'h c3ed80;
		246: head_rom_data = 24'h c3ed80;
		247: head_rom_data = 24'h c3ed80;
		248: head_rom_data = 24'h c3ed80;
		249: head_rom_data = 24'h c3ed80;
		250: head_rom_data = 24'h c3ed80;
		251: head_rom_data = 24'h c3ed80;
		252: head_rom_data = 24'h 074b2b;
		253: head_rom_data = 24'h 1a1a1c;
		254: head_rom_data = 24'h 1a1a1c;
		255: head_rom_data = 24'h 1a1a1c;
		default: ;
	endcase
end

endmodule